module multiply_sim(

    );
endmodule